------------------------------------------------------------------------------
-- Noridel Herron
-- 7/16/2025
-- MEM_WB Register
------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use IEEE.MATH_REAL.ALL;

-- CUSTOM PACKAGES
library work;
use work.Pipeline_Types.all;
use work.const_Types.all;
use work.initialize_records.all;
use work.ENUM_T.all;
--use work.MyFunctions.all;
entity MEM_WB is
    Port ( 
           clk            : in   std_logic; 
           reset          : in   std_logic;
           -- inputs from ex_mem register
           ex_mem         : in  Inst_PC_N;
           exmem_content  : in  EX_CONTENT_N;
           -- inputs from mem stage
           memA_result    : in  std_logic_vector(DATA_WIDTH-1 downto 0); 
           -- outputs
           mem_wb         : out Inst_PC_N;  
           mem_wb_content : out MEM_CONTENT_N  
        );
        
end MEM_WB;

architecture Behavioral of MEM_WB is

signal reg         : Inst_PC_N      := EMPTY_Inst_PC_N;
signal reg_content : MEM_CONTENT_N  := EMPTY_MEM_CONTENT_N;

begin
    process(clk, reset)
    variable reg_content_v : MEM_CONTENT_N := EMPTY_MEM_CONTENT_N;
    begin
        if reset = '1' then  
            -- clear everything
            reg         <= EMPTY_Inst_PC_N;
            reg_content <= EMPTY_MEM_CONTENT_N;
        
        elsif rising_edge(clk) then
            reg               <= ex_mem;
            -- A contents
            reg_content_v.A.alu := exmem_content.A.alu.result;
            reg_content_v.A.rd  := exmem_content.A.rd;
            reg_content_v.A.we  := exmem_content.A.cntrl.wb;
            reg_content_v.A.me  := exmem_content.A.cntrl.mem;
            reg_content_v.A.mem := (others => '0');
            
            -- B contents 
            reg_content_v.B.alu := exmem_content.B.alu.result;
            reg_content_v.B.rd  := exmem_content.B.rd;
            reg_content_v.B.we  := exmem_content.B.cntrl.wb;
            reg_content_v.B.me  := exmem_content.B.cntrl.mem;
            reg_content_v.B.mem := (others => '0');
            
            if ex_mem.isMemBusy = MEM_A and (exmem_content.A.cntrl.mem = MEM_READ or exmem_content.A.cntrl.mem = MEM_WRITE) then
                reg_content_v.A.mem := memA_result;
            
            elsif ex_mem.isMemBusy = MEM_B and (exmem_content.B.cntrl.mem = MEM_READ or exmem_content.B.cntrl.mem = MEM_WRITE) then
                reg_content_v.B.mem := memA_result;
            
            elsif (exmem_content.A.cntrl.mem = MEM_READ or exmem_content.A.cntrl.mem = MEM_WRITE) then
                reg_content_v.A.mem := memA_result;
                
            elsif (exmem_content.B.cntrl.mem = MEM_READ or exmem_content.B.cntrl.mem = MEM_WRITE) then
                reg_content_v.B.mem := memA_result;  
            end if;
            reg_content <= reg_content_v;
        end if;    
    end process;

    -- assign output
    mem_wb         <= reg;
    mem_wb_content <= reg_content;

end Behavioral;