`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 06/18/2025 10:13:07 AM
// Design Name: Noridel Herron
// Module Name: EX_STAGE
// Project Name: Superscalar CPU
//////////////////////////////////////////////////////////////////////////////////


module EX_STAGE(

    );
endmodule
